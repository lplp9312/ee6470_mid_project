`timescale 1ps / 1ps
/*****************************************************************************
    Verilog RTL Description
    
    Configured at: 00:40:24 CST (+0800), Wednesday 05 May 2021
    Configured on: ws28
    Configured by: m109061634 (m109061634)
    
    Created by: Stratus DpOpt 2019.1.01 
*******************************************************************************/

module DC_Filter_gen000002_4 (
	in1,
	out1
	); /* architecture "behavioural" */ 
input [8:0] in1;
output [10:0] out1;
wire [10:0] asc001;

assign asc001 = 
	+(in1)
	+(11'B01000000100);

assign out1 = asc001;
endmodule

/* CADENCE  ubHzQgs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE ******/


